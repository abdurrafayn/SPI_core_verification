package spi_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "spi_packet.sv"
    `include "spi_driver.sv"
    `include "spi_monitor.sv"
    `include "spi_sequencer.sv"
    `include "spi_agent.sv"
    `include "spi_env.sv"


endpackage