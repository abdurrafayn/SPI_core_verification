package wb_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "wb_packet.sv"
    `include "wb_driver.sv"
    `include "wb_monitor.sv"
    `include "wb_sequencer.sv"
    `include "wb_agent.sv"


endpackage